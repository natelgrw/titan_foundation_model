.suckt  two_stage_fully_differential_op_amp_23_3 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
mDiodeTransistorPmos3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mDiodeTransistorPmos4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos8 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos9 out1 out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos10 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos11 out2 out2FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos12 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos13 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos15 sourceTransconductance ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos16 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos17 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos18 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos19 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos20 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos21 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
mNormalTransistorPmos22 out1 inputVoltageBiasXXpXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
mNormalTransistorPmos23 out1FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mNormalTransistorPmos24 out2 inputVoltageBiasXXpXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
mNormalTransistorPmos25 out2FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos26 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos27 FirstStageYinnerTransistorStack1Load2 outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos28 FirstStageYinnerTransistorStack2Load2 outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos29 SecondStage1YinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos30 SecondStage2YinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_23_3

