.suckt  two_stage_single_output_op_amp_67_10 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorPmos3 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mDiodeTransistorPmos6 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 FirstStageYinnerOutputLoad2 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos11 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos12 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorPmos13 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mNormalTransistorPmos14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos15 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos16 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos17 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos18 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos
mNormalTransistorPmos19 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos20 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos21 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
mNormalTransistorPmos22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_67_10

