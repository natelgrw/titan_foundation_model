.suckt  one_stage_fully_differential_op_amp63 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorPmos5 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos8 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos9 out1 outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
mNormalTransistorNmos10 out2 outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mNormalTransistorNmos11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos15 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos16 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos17 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos18 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos19 FirstStageYinnerTransistorStack1Load2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos20 FirstStageYinnerTransistorStack2Load2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos21 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos22 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos23 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos24 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos25 out1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mNormalTransistorPmos26 out2 outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mNormalTransistorPmos27 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos28 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos29 FirstStageYsourceGCC1 outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos30 FirstStageYsourceGCC2 outFeedback sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out2 sourceNmos 
.end one_stage_fully_differential_op_amp63

