.suckt  one_stage_fully_differential_op_amp44 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos
mDiodeTransistorPmos5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mDiodeTransistorPmos6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mDiodeTransistorPmos8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos
mNormalTransistorNmos9 out1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos10 out2 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos11 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos12 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorPmos13 out1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mNormalTransistorPmos14 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorPmos15 out2 outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mNormalTransistorPmos16 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos17 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos18 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mNormalTransistorPmos19 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorPmos20 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorPmos21 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos22 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos23 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
mNormalTransistorPmos24 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
mNormalTransistorPmos25 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos26 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos27 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out2 sourceNmos 
.end one_stage_fully_differential_op_amp44

