.suckt  two_stage_single_output_op_amp_127_7 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos2 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos4 out inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos5 outFirstStage inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos6 FirstStageYout1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos7 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos8 out outFirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos9 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorPmos10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_127_7

