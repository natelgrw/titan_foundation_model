.suckt  one_stage_fully_differential_op_amp69 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
mDiodeTransistorPmos4 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos8 out1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos9 out2 outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos12 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos14 sourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
mNormalTransistorNmos15 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos16 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos17 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos18 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos19 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos20 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos21 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
mNormalTransistorPmos22 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos23 out1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mNormalTransistorPmos24 out2 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos25 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos26 FirstStageYinnerTransistorStack1Load2 outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos27 FirstStageYinnerTransistorStack2Load2 outFeedback sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out2 sourceNmos 
.end one_stage_fully_differential_op_amp69

