.suckt  symmetrical_op_amp197 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mDiodeTransistorNmos3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mDiodeTransistorPmos5 out1FirstStage out1FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mNormalTransistorNmos6 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos7 out innerComplementarySecondStage sourceNmos sourceNmos nmos
mNormalTransistorNmos8 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
mNormalTransistorPmos11 innerComplementarySecondStage inSourceTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
mNormalTransistorPmos12 out out1FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mNormalTransistorPmos13 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos14 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mNormalTransistorPmos15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
.end symmetrical_op_amp197

