************************************************************************
* auCdl Netlist:
* 
* Library Name:  OTA_class
* Top Cell Name: fully_differential_gain_boosting
* View Name:     schematic
* Netlisted on:  Sep 11 21:05:36 2019
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!
+        gnd!

*.PIN vdd!
*+    gnd!

************************************************************************
* Library Name: OTA_class
* Cell Name:    fully_differential
* View Name:    schematic
************************************************************************

.SUBCKT fully_differential Vinn Vinp Voutn Voutp
*.PININFO Vinn:I Vinp:I Voutn:O Voutp:O
MM1 Voutn Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA1
MM2 Voutp Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA1
MM4 net14 Vbiasn gnd! gnd! nmos w=WA l=LA nfin=nA2
MM3 Voutn Vinp net14 gnd! nmos w=WA l=LA nfin=nA3
MM0 Voutp Vinn net14 gnd! nmos w=WA l=LA nfin=nA3
.ENDS

************************************************************************
* Library Name: OTA_class
* Cell Name:    fully_differential_gain_boosting
* View Name:    schematic
************************************************************************

.SUBCKT fully_differential_gain_boosting Vbiasn Vbiasp Vinn Vinp Voutn Voutp
*.PININFO Vbiasn:I Vbiasp:O Vinn:I Vinp:I Voutn:O Voutp:O
MM8 Voutn net22 net23 gnd! nmos w=WA l=LA nfin=nA1
MM7 Voutp net19 net21 gnd! nmos w=WA l=LA nfin=nA1
MM3 net23 Vinp net15 gnd! nmos w=WA l=LA nfin=nA2
MM0 net21 Vinn net15 gnd! nmos w=WA l=LA nfin=nA2
MM4 net15 Vbiasn gnd! gnd! nmos w=WA l=LA nfin=nA3
MM6 Voutn net24 net25 vdd pmos w=WA l=LA nfin=nA4
MM5 Voutp net20 net12 vdd pmos w=WA l=LA nfin=nA4
MM1 net25 Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA5
MM2 net12 Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA5
XI3 net12 net25 net24 net20 / fully_differential
XI1 net23 net21 net19 net22 / fully_differential
.ENDS


.SUBCKT LG_npmos Biasn Vbiasn Vbiasp
*.PININFO Biasn:I Vbiasn:O Vbiasp:O
MM4 Vbiasp Vbiasn gnd! gnd! nmos w=WA l=LA nfin=nA1
MM2 Vbiasn Vbiasn gnd! gnd! nmos w=WA l=LA nfin=nA2
MM10 neta Biasn gnd! gnd! nmos w=WA l=LA nfin=nA3
MM3 Vbiasp Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA4
MM1 Vbiasn neta vdd! vdd! pmos w=WA l=LA nfin=nA5
MM0 neta neta vdd! vdd! pmos w=WA l=LA nfin=nA5
.ENDS

.SUBCKT CR11_1 Vbiasn
*.PININFO Vbiasn:O
RRF vdd! Vbiasn res=rK
MM1 net9 Vbiasn gnd! gnd! nmos w=WA l=LA nfin=nA1
MM0 Vbiasn Vbiasn gnd! gnd! nmos w=WA l=LA nfin=nA1
MM3 net9 net9 vdd! vdd! pmos w=WA l=LA nfin=nA2
MM2 Vbiasn net9 vdd! vdd! pmos w=WA l=LA nfin=nA2
.ENDS


xiota LG_Vbiasn LG_Vbiasp Vinn Vinp Voutn Voutp fully_differential_gain_boosting
xiLG_npmos Biasn LG_Vbiasn LG_Vbiasp LG_npmos
xibCR11_1 Biasn CR11_1
.END