.suckt  two_stage_fully_differential_op_amp_14_11 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos3 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos4 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos8 out1 outVoltageBiasXXnXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias nmos
mNormalTransistorNmos9 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos10 out2 outVoltageBiasXXnXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias nmos
mNormalTransistorNmos11 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos15 FeedbackStageYinnerStageBias2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos16 FeedbackStageYinnerStageBias1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos17 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos18 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos19 FeedbackStageYsourceTransconductance1 outVoltageBiasXXnXX1 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
mNormalTransistorNmos20 FeedbackStageYsourceTransconductance2 outVoltageBiasXXnXX1 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
mNormalTransistorNmos21 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos22 SecondStage1YinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos23 SecondStage2YinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorPmos24 out1 outVoltageBiasXXpXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
mNormalTransistorPmos25 out1FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos26 out2 outVoltageBiasXXpXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
mNormalTransistorPmos27 out2FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos28 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos29 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos30 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_14_11

