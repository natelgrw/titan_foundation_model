.suckt  two_stage_single_output_op_amp_86_3 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos
mDiodeTransistorPmos3 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorNmos6 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos7 out outFirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos
mNormalTransistorNmos9 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos
mNormalTransistorPmos11 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos12 out outVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mNormalTransistorPmos13 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mNormalTransistorPmos14 sourceTransconductance ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mNormalTransistorPmos16 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos17 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos18 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_86_3

