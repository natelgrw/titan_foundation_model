.suckt  complementary_op_amp15 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorPmos3 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorNmos5 out inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
mNormalTransistorNmos6 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos7 FirstStageYinnerStageBiasNmos outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos8 FirstStageYinnerTransistorStack1LoadNmos FirstStageYout1 sourceNmos sourceNmos nmos
mNormalTransistorNmos9 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
mNormalTransistorNmos10 FirstStageYinnerTransistorStack2LoadNmos FirstStageYout1 sourceNmos sourceNmos nmos
mNormalTransistorNmos11 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
mNormalTransistorNmos12 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
mNormalTransistorNmos13 FirstStageYsourceTransconductanceNmos inputVoltageBiasXXnXX1 FirstStageYinnerStageBiasNmos FirstStageYinnerStageBiasNmos nmos
mNormalTransistorPmos14 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
mNormalTransistorPmos15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos16 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos17 FirstStageYinnerStageBiasPmos ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos18 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
mNormalTransistorPmos19 FirstStageYinnerTransistorStack1LoadPmos FirstStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorPmos20 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
mNormalTransistorPmos21 FirstStageYinnerTransistorStack2LoadPmos FirstStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorPmos22 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
mNormalTransistorPmos23 FirstStageYsourceTransconductancePmos outVoltageBiasXXpXX1 FirstStageYinnerStageBiasPmos FirstStageYinnerStageBiasPmos pmos
Capacitor1 out sourceNmos 
.end complementary_op_amp15

