.suckt  one_stage_single_output_op_amp1 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos2 ibias ibias sourcePmos sourcePmos pmos
mNormalTransistorNmos3 out FirstStageYout1 sourceNmos sourceNmos nmos
mNormalTransistorPmos4 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos6 out in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
Capacitor1 out sourceNmos 
.end one_stage_single_output_op_amp1

