.suckt  two_stage_fully_differential_op_amp_24_9 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX4 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
mDiodeTransistorNmos5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos7 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos
mDiodeTransistorPmos8 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos9 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos10 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos11 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos12 out1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos13 out1FirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos14 out2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
mNormalTransistorNmos15 out2FirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos16 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos17 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos18 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos19 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos20 sourceTransconductance ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos21 FeedbackStageYinnerStageBias1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos22 FeedbackStageYinnerStageBias2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos23 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos24 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos25 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX4 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
mNormalTransistorNmos26 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX4 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
mNormalTransistorNmos27 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos28 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos29 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos30 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorPmos31 inputVoltageBiasXXnXX4 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos32 out1 out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos33 out1FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mNormalTransistorPmos34 out2 out2FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos35 out2FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos36 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos37 outInputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos38 outVoltageBiasXXnXX3 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos39 FirstStageYinnerTransistorStack1Load2 outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos40 FirstStageYinnerTransistorStack2Load2 outFeedback sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_24_9

