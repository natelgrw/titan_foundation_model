************************************************************************
* auCdl Netlist:
* 
* Library Name:  OTA_class
* Top Cell Name: single_ended_low_voltage_cascode_pmos
* View Name:     schematic
* Netlisted on:  Sep 11 21:08:22 2019
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!
+        gnd!

*.PIN vdd!
*+    gnd!

************************************************************************
* Library Name: OTA_class
* Cell Name:    single_ended_low_voltage_cascode_pmos
* View Name:    schematic
************************************************************************

.SUBCKT single_ended_low_voltage_cascode_pmos Vbiasp Vinn Vinp Voutp
*.PININFO Vbiasp:I Vinn:I Vinp:I Voutp:O
MM7 Voutp Vinn net11 net18 pmos w=WA l=LA nfin=nA1
MM6 net13 Vinp net11 net18 pmos w=WA l=LA nfin=nA1
MM5 net11 Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA2
MM1 Voutp net17 net20 gnd! nmos w=WA l=LA nfin=nA3
MM0 net13 net17 net19 gnd! nmos w=WA l=LA nfin=nA3
MM9 net20 net13 gnd! gnd! nmos w=WA l=LA nfin=nA4
MM8 net19 net13 gnd! gnd! nmos w=WA l=LA nfin=nA4
.ENDS


.SUBCKT LG_pmos Biasn Vbiasp
*.PININFO Biasn:I Vbiasp:O
MM10 Vbiasp Biasn gnd! gnd! nmos w=WA l=LA nfin=nA1
MM3 Vbiasp Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA2
.ENDS

.SUBCKT CR12_1 Vbiasn
*.PININFO Vbiasn:O
MM0 Vbiasn Vbiasn gnd! gnd! nmos w=WA l=LA nfin=nA1
MM1 net10 Vbiasn gnd! gnd! nmos w=WA l=LA nfin=nA1
MM2 Vbiasn net10 vdd! vdd! pmos w=WA l=LA nfin=nA2
RRF vdd! Vbiasn res=rK
RR0 vdd! net10 res=rK
.ENDS


xiota LG_Vbiasp Vinn Vinp Voutp single_ended_low_voltage_cascode_pmos
xiLG_pmos Biasn LG_Vbiasp LG_pmos
xibCR12_1 Biasn CR12_1
.END