.suckt  two_stage_fully_differential_op_amp_42_10 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
mDiodeTransistorPmos6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 out1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos8 inputVoltageBiasXXpXX3 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos9 out1FirstStage outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos10 out2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos11 out2FirstStage outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos13 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mNormalTransistorPmos14 out1 outVoltageBiasXXpXX2 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
mNormalTransistorPmos15 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mNormalTransistorPmos16 out2 outVoltageBiasXXpXX2 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
mNormalTransistorPmos17 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mNormalTransistorPmos18 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos19 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos20 sourceTransconductance outVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
mNormalTransistorPmos21 FeedbackStageYinnerStageBias2 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorPmos22 FeedbackStageYinnerStageBias1 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorPmos23 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos24 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos25 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
mNormalTransistorPmos26 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
mNormalTransistorPmos27 FirstStageYinnerStageBias inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorPmos28 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos29 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos30 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos31 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_42_10

