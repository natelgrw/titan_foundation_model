.suckt  two_stage_fully_differential_op_amp_32_11 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mDiodeTransistorPmos6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mDiodeTransistorPmos8 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorNmos9 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias nmos
mNormalTransistorNmos10 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mNormalTransistorNmos11 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias nmos
mNormalTransistorNmos12 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mNormalTransistorNmos13 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos15 outVoltageBiasXXpXX3 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos16 FirstStageYinnerTransistorStack1Load1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos17 FirstStageYinnerTransistorStack2Load1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos18 SecondStage1YinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos19 SecondStage2YinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorPmos20 out1 outVoltageBiasXXpXX2 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
mNormalTransistorPmos21 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorPmos22 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos23 out2 outVoltageBiasXXpXX2 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
mNormalTransistorPmos24 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos25 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos26 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos27 FeedbackStageYinnerStageBias1 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorPmos28 FeedbackStageYinnerStageBias2 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mNormalTransistorPmos29 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos30 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos31 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
mNormalTransistorPmos32 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
mNormalTransistorPmos33 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mNormalTransistorPmos34 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos35 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos36 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_32_11

