.suckt  two_stage_fully_differential_op_amp_12_1 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos5 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
mNormalTransistorNmos8 inputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos9 out1 out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos10 out1FirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
mNormalTransistorNmos11 out2 out2FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos12 out2FirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mNormalTransistorNmos13 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos14 FirstStageYinnerTransistorStack1Load2 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos15 FirstStageYinnerTransistorStack2Load2 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorPmos16 out1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos17 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mNormalTransistorPmos18 out2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos19 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mNormalTransistorPmos20 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos21 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos22 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos23 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos24 sourceTransconductance ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos25 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos26 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos27 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos28 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos29 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXpXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
mNormalTransistorPmos30 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXpXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
mNormalTransistorPmos31 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos32 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_12_1

