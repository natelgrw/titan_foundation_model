.suckt  two_stage_fully_differential_op_amp_47_2 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos5 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos
mDiodeTransistorPmos7 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mDiodeTransistorPmos8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorNmos9 inputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
mNormalTransistorNmos11 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
mNormalTransistorNmos12 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
mNormalTransistorNmos13 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mNormalTransistorNmos14 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos15 FirstStageYinnerTransistorStack1Load2 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos16 FirstStageYinnerTransistorStack2Load2 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos17 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos18 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
mNormalTransistorPmos19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos20 out1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos21 out1FirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mNormalTransistorPmos22 out2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos23 out2FirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mNormalTransistorPmos24 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos25 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos26 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos27 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mNormalTransistorPmos28 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos29 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos30 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos31 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos32 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos33 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos34 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_47_2

