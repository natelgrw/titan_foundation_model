.suckt  two_stage_fully_differential_op_amp_71_3 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos
mDiodeTransistorPmos5 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos8 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos9 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 out1 out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos11 out1FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos12 out2 out2FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos13 out2FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos14 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos15 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos16 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos17 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos18 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos19 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mNormalTransistorNmos20 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mNormalTransistorNmos21 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos22 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos23 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos24 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos25 out1 inputVoltageBiasXXpXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
mNormalTransistorPmos26 out1FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mNormalTransistorPmos27 out2 inputVoltageBiasXXpXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
mNormalTransistorPmos28 out2FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos29 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos30 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos31 FirstStageYinnerTransistorStack1Load2 outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos32 FirstStageYinnerTransistorStack2Load2 outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos33 SecondStage1YinnerStageBias ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos34 SecondStage2YinnerStageBias ibias sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_71_3

