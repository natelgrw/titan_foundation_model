.suckt  symmetrical_op_amp89 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage nmos
mDiodeTransistorNmos2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 out1FirstStage out1FirstStage sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 out2FirstStage out2FirstStage out1FirstStage out1FirstStage nmos
mDiodeTransistorPmos5 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
mNormalTransistorNmos7 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
mNormalTransistorNmos8 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mNormalTransistorNmos9 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos10 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mNormalTransistorPmos11 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos12 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mNormalTransistorPmos13 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos15 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos
mNormalTransistorPmos16 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
.end symmetrical_op_amp89

