.suckt  two_stage_single_output_op_amp_34_6 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mDiodeTransistorPmos5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mDiodeTransistorPmos8 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 out inputVoltageBiasXXnXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mNormalTransistorNmos11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos12 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos14 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos15 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos16 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos17 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos18 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos19 out inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mNormalTransistorPmos20 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mNormalTransistorPmos21 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorPmos22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_34_6

