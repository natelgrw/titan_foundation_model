.suckt  two_stage_fully_differential_op_amp_66_10 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
mDiodeTransistorPmos4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos8 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos9 out1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos10 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos11 out2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos12 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos13 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos16 sourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
mNormalTransistorNmos17 FeedbackStageYinnerStageBias1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos18 FeedbackStageYinnerStageBias2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos19 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos20 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos21 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
mNormalTransistorNmos22 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
mNormalTransistorNmos23 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos24 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos25 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
mNormalTransistorPmos26 inputVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos27 out1 outVoltageBiasXXpXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
mNormalTransistorPmos28 out1FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos29 out2 outVoltageBiasXXpXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
mNormalTransistorPmos30 out2FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos31 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos32 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos33 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_66_10

