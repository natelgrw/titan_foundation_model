.suckt  two_stage_single_output_op_amp_97_9 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mNormalTransistorNmos8 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos9 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos11 sourceTransconductance ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos12 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos
mNormalTransistorPmos17 out outFirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos18 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos19 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos20 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos
Capacitor1 outFirstStage out 
Capacitor2 out sourceNmos 
.end two_stage_single_output_op_amp_97_9

