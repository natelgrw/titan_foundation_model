.suckt  two_stage_fully_differential_op_amp_49_2 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorPmos3 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos4 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos6 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
mNormalTransistorNmos7 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos8 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
mNormalTransistorNmos9 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos12 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos14 FeedbackStageYsourceTransconductance1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos15 FeedbackStageYsourceTransconductance2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos16 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos17 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
mNormalTransistorNmos18 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos19 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
mNormalTransistorPmos20 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos21 out1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos22 out1FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos23 out2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos24 out2FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos25 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_49_2

