.suckt  two_stage_single_output_op_amp_146_2 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorNmos6 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mNormalTransistorNmos7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mNormalTransistorNmos8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos9 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos10 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos11 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourceNmos sourceNmos nmos
mNormalTransistorNmos12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos13 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos14 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
mNormalTransistorPmos15 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos16 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos17 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos18 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos19 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos20 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_146_2

