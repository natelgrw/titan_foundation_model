.suckt  two_stage_fully_differential_op_amp_40_9 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
mDiodeTransistorNmos4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos6 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos7 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mDiodeTransistorNmos8 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos9 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
mDiodeTransistorPmos10 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mDiodeTransistorPmos11 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos12 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorNmos13 out1FirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos14 out1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos15 out2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
mNormalTransistorNmos16 out2FirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos17 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos18 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos19 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos20 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos21 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorPmos22 out1FirstStage ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mNormalTransistorPmos23 out1 out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos24 out2 out2FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos25 out2FirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos26 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos27 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos28 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos29 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos30 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos31 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos32 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos33 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos34 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos35 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos36 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
mNormalTransistorPmos37 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
mNormalTransistorPmos38 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos39 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos40 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos41 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos42 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mNormalTransistorPmos43 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
Capacitor1 out1FirstStage out1 
Capacitor2 out1 sourceNmos 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_40_9

