.suckt  two_stage_fully_differential_op_amp_4_5 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos5 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mDiodeTransistorPmos7 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mDiodeTransistorPmos8 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
mDiodeTransistorPmos9 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos10 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorNmos11 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos12 inputVoltageBiasXXpXX3 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos13 out1 out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos14 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mNormalTransistorNmos15 out2 out2FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos16 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mNormalTransistorNmos17 outInputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos18 FirstStageYinnerTransistorStack1Load1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos19 FirstStageYinnerTransistorStack2Load1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorPmos20 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos21 out1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mNormalTransistorPmos22 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos23 out2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
mNormalTransistorPmos24 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos25 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos26 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos27 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos28 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos29 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos30 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos31 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos32 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXpXX3 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
mNormalTransistorPmos33 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXpXX3 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
mNormalTransistorPmos34 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos35 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorPmos36 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_4_5

