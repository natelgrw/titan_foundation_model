.suckt  two_stage_fully_differential_op_amp_42_1 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
mNormalTransistorNmos7 out1 out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos8 out2 out2FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos9 out1FirstStage outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos10 inputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos11 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos12 out2FirstStage outFeedback sourceNmos sourceNmos nmos
mNormalTransistorPmos13 out1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos14 out2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos15 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mNormalTransistorPmos16 sourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
mNormalTransistorPmos17 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos18 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos19 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos20 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mNormalTransistorPmos21 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos22 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos23 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos24 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos25 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXpXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
mNormalTransistorPmos26 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXpXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
mNormalTransistorPmos27 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos28 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
mNormalTransistorPmos29 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out2 sourceNmos 
Capacitor3 out1FirstStage out1 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_42_1

