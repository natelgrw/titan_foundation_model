.suckt  two_stage_single_output_op_amp_205_2 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mDiodeTransistorPmos5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos8 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos9 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mNormalTransistorNmos10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos
mNormalTransistorNmos11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos12 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos13 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos
mNormalTransistorNmos14 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos15 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
mNormalTransistorNmos16 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
mNormalTransistorPmos17 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos18 out inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos20 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos21 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos22 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_205_2

