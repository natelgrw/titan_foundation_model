.suckt  symmetrical_op_amp92 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos
mDiodeTransistorPmos2 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos3 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos
mNormalTransistorNmos4 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mNormalTransistorNmos5 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
mNormalTransistorNmos6 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mNormalTransistorNmos7 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mNormalTransistorNmos8 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos9 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mNormalTransistorNmos10 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos11 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mNormalTransistorPmos12 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos13 out innerComplementarySecondStage sourcePmos sourcePmos pmos
mNormalTransistorPmos14 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos15 out2FirstStage ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
.end symmetrical_op_amp92

