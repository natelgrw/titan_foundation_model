.suckt  two_stage_single_output_op_amp_141_5 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 FirstStageYinnerLoad1 FirstStageYinnerLoad1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mDiodeTransistorPmos4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorNmos6 out outFirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos7 outFirstStage FirstStageYinnerLoad1 sourceNmos sourceNmos nmos
mNormalTransistorNmos8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos9 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos10 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos11 FirstStageYinnerLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos12 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mNormalTransistorPmos13 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mNormalTransistorPmos14 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos15 FirstStageYinnerLoad1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mNormalTransistorPmos16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_141_5

