.suckt  two_stage_fully_differential_op_amp_14_1 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorPmos3 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos4 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos6 out1 out1FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos7 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos8 out2 out2FirstStage sourceNmos sourceNmos nmos
mNormalTransistorNmos9 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos12 FeedbackStageYinnerStageBias1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos13 FeedbackStageYinnerStageBias2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos14 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos15 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos16 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX1 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
mNormalTransistorNmos17 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX1 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
mNormalTransistorNmos18 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorPmos19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos20 out1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos21 out1FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos22 out2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos23 out2FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos24 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_14_1

