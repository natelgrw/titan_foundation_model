.suckt  two_stage_fully_differential_op_amp_68_7 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos
mDiodeTransistorPmos6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos7 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos8 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos10 out1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos11 out1FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos12 out2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos13 out2FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos14 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos15 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos16 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos17 FeedbackStageYinnerStageBias1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos18 FeedbackStageYinnerStageBias2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos19 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos20 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos21 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX3 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
mNormalTransistorNmos22 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX3 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
mNormalTransistorNmos23 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos24 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos25 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos26 inputVoltageBiasXXnXX3 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos27 out1 out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos28 out1FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos29 out2 out2FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos30 out2FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos31 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos32 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_68_7

