.suckt  two_stage_fully_differential_op_amp_21_8 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 out1 outVoltageBiasXXnXX2 SecondStage1YinnerStageBias SecondStage1YinnerStageBias nmos
mNormalTransistorNmos8 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos9 out2 outVoltageBiasXXnXX2 SecondStage2YinnerStageBias SecondStage2YinnerStageBias nmos
mNormalTransistorNmos10 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos14 sourceTransconductance ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos15 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos16 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos17 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos18 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos19 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos20 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos21 SecondStage1YinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos22 SecondStage2YinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorPmos23 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos24 out1 out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos25 out1FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos26 out2 out2FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos27 out2FirstStage outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos28 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_21_8

