.suckt  two_stage_single_output_op_amp_139_1 outVoltageBiasXXpXX1 in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos2 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mDiodeTransistorPmos3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorNmos4 FirstStageYinnerOutputLoad1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos5 outFirstStage outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos6 out outFirstStage sourceNmos sourceNmos nmos
mNormalTransistorPmos7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerOutputLoad1 sourcePmos sourcePmos pmos
mNormalTransistorPmos8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerOutputLoad1 sourcePmos sourcePmos pmos
mNormalTransistorPmos10 outVoltageBiasXXnXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorPmos11 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mNormalTransistorPmos12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos13 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorPmos14 out outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
Capacitor1 outFirstStage out 
Capacitor2 out sourceNmos 
.end two_stage_single_output_op_amp_139_1

