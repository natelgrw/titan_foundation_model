.suckt  symmetrical_op_amp200 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorPmos3 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mDiodeTransistorPmos4 out1FirstStage out1FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorNmos6 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos7 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos
mNormalTransistorNmos8 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
mNormalTransistorNmos9 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos11 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos12 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
mNormalTransistorNmos13 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
mNormalTransistorNmos14 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos
mNormalTransistorPmos15 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos16 innerComplementarySecondStage inSourceTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
mNormalTransistorPmos17 out out1FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mNormalTransistorPmos18 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos19 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mNormalTransistorPmos20 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos21 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
.end symmetrical_op_amp200

