.suckt  one_stage_single_output_op_amp127 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos2 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos3 ibias ibias sourcePmos sourcePmos pmos
mNormalTransistorNmos4 FirstStageYout1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos5 out outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos6 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos8 out in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos9 out FirstStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorPmos10 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
.end one_stage_single_output_op_amp127

