.suckt  complementary_op_amp29 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mDiodeTransistorNmos2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 FirstStageYinnerOutputLoadNmos FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
mDiodeTransistorNmos4 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos sourceNmos sourceNmos nmos
mDiodeTransistorPmos5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mDiodeTransistorPmos6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 out FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
mNormalTransistorNmos8 FirstStageYinnerStageBiasNmos outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos9 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
mNormalTransistorNmos10 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack1LoadNmos sourceNmos sourceNmos nmos
mNormalTransistorNmos11 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
mNormalTransistorNmos12 FirstStageYsourceTransconductanceNmos outInputVoltageBiasXXnXX1 FirstStageYinnerStageBiasNmos FirstStageYinnerStageBiasNmos nmos
mNormalTransistorPmos13 out ibias FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
mNormalTransistorPmos14 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorPmos15 FirstStageYinnerOutputLoadNmos ibias FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
mNormalTransistorPmos16 FirstStageYinnerStageBiasPmos outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorPmos17 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
mNormalTransistorPmos18 FirstStageYinnerTransistorStack1LoadPmos outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorPmos19 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
mNormalTransistorPmos20 FirstStageYinnerTransistorStack2LoadPmos outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorPmos21 FirstStageYsourceTransconductancePmos ibias FirstStageYinnerStageBiasPmos FirstStageYinnerStageBiasPmos pmos
Capacitor1 out sourceNmos 
.end complementary_op_amp29

