.suckt  two_stage_single_output_op_amp_129_12 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos8 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos9 outFirstStage outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 FirstStageYout1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos12 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mNormalTransistorPmos13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos
mNormalTransistorPmos14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos15 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos16 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos17 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mNormalTransistorPmos18 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos19 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_129_12

