.suckt  two_stage_fully_differential_op_amp_29_9 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos3 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
mDiodeTransistorNmos5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos7 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos8 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos9 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos10 ibias ibias sourcePmos sourcePmos pmos
mNormalTransistorNmos11 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos12 out1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos13 out1FirstStage inputVoltageBiasXXnXX3 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mNormalTransistorNmos14 out2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
mNormalTransistorNmos15 out2FirstStage inputVoltageBiasXXnXX3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mNormalTransistorNmos16 FirstStageYinnerTransistorStack1Load1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos17 FirstStageYinnerTransistorStack2Load1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos18 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos19 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorPmos20 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos21 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos22 out1 out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos23 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos24 out2 out2FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos25 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos26 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos27 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos28 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos29 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos30 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos31 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos32 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos33 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos34 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos35 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_29_9

