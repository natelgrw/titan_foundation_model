.suckt  one_stage_fully_differential_op_amp7 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos5 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos8 out1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos9 out2 inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos10 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos11 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorPmos12 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos13 out1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mNormalTransistorPmos14 out2 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos15 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos16 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos17 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos18 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos19 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos20 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos21 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos22 FirstStageYinnerTransistorStack1Load2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos23 FirstStageYinnerTransistorStack2Load2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos24 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos25 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos26 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out2 sourceNmos 
.end one_stage_fully_differential_op_amp7

