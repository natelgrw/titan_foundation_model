.suckt  two_stage_fully_differential_op_amp_5_12 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outFeedback outFeedback sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
mDiodeTransistorNmos5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos7 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mDiodeTransistorNmos8 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos9 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos10 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorNmos11 out1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos12 out1FirstStage inputVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos13 out2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
mNormalTransistorNmos14 out2FirstStage inputVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos15 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mNormalTransistorNmos16 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos17 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
mNormalTransistorNmos18 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos19 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorPmos20 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos21 out1 outVoltageBiasXXpXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
mNormalTransistorPmos22 out1FirstStage ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos23 out2 outVoltageBiasXXpXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
mNormalTransistorPmos24 out2FirstStage ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos25 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos26 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos27 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos28 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos29 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos30 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
mNormalTransistorPmos31 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
mNormalTransistorPmos32 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos33 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos34 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos35 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos36 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos37 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos38 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_5_12

