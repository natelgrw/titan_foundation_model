.suckt  complementary_op_amp10 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorPmos3 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorNmos5 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos6 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
mNormalTransistorNmos7 FirstStageYinnerSourceLoadNmos outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
mNormalTransistorNmos8 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
mNormalTransistorNmos9 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
mNormalTransistorNmos10 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
mNormalTransistorNmos11 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
mNormalTransistorNmos12 FirstStageYsourceTransconductanceNmos inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorPmos13 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos14 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
mNormalTransistorPmos15 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos16 FirstStageYinnerSourceLoadNmos inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
mNormalTransistorPmos17 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
mNormalTransistorPmos18 FirstStageYinnerTransistorStack1LoadPmos ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos19 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
mNormalTransistorPmos20 FirstStageYinnerTransistorStack2LoadPmos ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos21 FirstStageYsourceTransconductancePmos ibias sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
.end complementary_op_amp10

