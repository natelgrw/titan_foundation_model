.suckt  two_stage_fully_differential_op_amp_19_12 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
mDiodeTransistorNmos1 ibias ibias sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
mDiodeTransistorNmos4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos6 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mDiodeTransistorPmos7 outFeedback outFeedback sourcePmos sourcePmos pmos
mDiodeTransistorPmos8 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mDiodeTransistorPmos9 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos10 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos11 out1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos12 out1FirstStage outVoltageBiasXXnXX3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
mNormalTransistorNmos13 out2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
mNormalTransistorNmos14 out2FirstStage outVoltageBiasXXnXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mNormalTransistorNmos15 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos16 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos17 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos18 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos19 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
mNormalTransistorNmos20 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
mNormalTransistorNmos21 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos22 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos23 FirstStageYinnerTransistorStack1Load2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos24 FirstStageYinnerTransistorStack2Load2 ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos25 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos26 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mNormalTransistorNmos27 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mNormalTransistorNmos28 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorNmos29 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorPmos30 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos31 out1 outVoltageBiasXXpXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
mNormalTransistorPmos32 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mNormalTransistorPmos33 out2 outVoltageBiasXXpXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
mNormalTransistorPmos34 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mNormalTransistorPmos35 outInputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos36 outVoltageBiasXXnXX3 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mNormalTransistorPmos37 FirstStageYsourceGCC1 outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos38 FirstStageYsourceGCC2 outFeedback sourcePmos sourcePmos pmos
mNormalTransistorPmos39 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos40 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
Capacitor1 out1 sourceNmos 
Capacitor2 out1FirstStage out1 
Capacitor3 out2 sourceNmos 
Capacitor4 out2FirstStage out2 
.end two_stage_fully_differential_op_amp_19_12

