.suckt  two_stage_single_output_op_amp_27_9 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mDiodeTransistorPmos4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mDiodeTransistorPmos5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorNmos6 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mNormalTransistorNmos7 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos8 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourceNmos sourceNmos nmos
mNormalTransistorNmos9 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos12 out outFirstStage sourcePmos sourcePmos pmos
mNormalTransistorPmos13 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorPmos14 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mNormalTransistorPmos15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos16 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
Capacitor1 outFirstStage out 
Capacitor2 out sourceNmos 
.end two_stage_single_output_op_amp_27_9

