************************************************************************
* auCdl Netlist:
* 
* Library Name:  OTA_class
* Top Cell Name: fully_differential_folded_cascode_pmos
* View Name:     schematic
* Netlisted on:  Sep 11 21:03:18 2019
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!
+        gnd!

*.PIN vdd!
*+    gnd!

************************************************************************
* Library Name: OTA_class
* Cell Name:    fully_differential_folded_cascode_pmos
* View Name:    schematic
************************************************************************

.SUBCKT fully_differential_folded_cascode_pmos Vbiasn1 Vbiasn2 Vbiasp Vbiasp1 Vbiasp2 Vinn Vinp Voutn Voutp
*.PININFO Vbiasn1:I Vbiasn2:I Vbiasp:I Vbiasp1:I Vbiasp2:I Vinn:I Vinp:I Voutn:O Voutp:O
MM8 Voutn Vbiasn2 net23 gnd! nmos w=WA l=LA nfin=nA1
MM7 Voutp Vbiasn2 net22 gnd! nmos w=WA l=LA nfin=nA1
MM10 net23 Vbiasn1 gnd! gnd! nmos w=WA l=LA nfin=nA2
MM9 net22 Vbiasn1 gnd! gnd! nmos w=WA l=LA nfin=nA2
MM0 net12 Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA3
MM2 net26 Vbiasp1 vdd! vdd! pmos w=WA l=LA nfin=nA4
MM1 net24 Vbiasp1 vdd! vdd! pmos w=WA l=LA nfin=nA4
MM4 net22 Vinn net12 net27 pmos w=WA l=LA nfin=nA5
MM3 net23 Vinp net12 net27 pmos w=WA l=LA nfin=nA5
MM6 Voutn Vbiasp2 net26 vdd! pmos w=WA l=LA nfin=nA6
MM5 Voutp Vbiasp2 net24 vdd! pmos w=WA l=LA nfin=nA6
.ENDS


.SUBCKT LG_load_biasn_LV Vbiasn2 Biasp
*.PININFO Vbiasn2:O Biasp:I 
MM13 net9 Vbiasn2 gnd! gnd! nmos w=WA l=LA nfin=nA1
MM15 Vbiasn2 Vbiasn2 net9 gnd! nmos w=WA l=LA nfin=nA2
MM14 Vbiasn2 Biasp vdd! vdd! pmos w=WA l=LA nfin=nA3
.ENDS

.SUBCKT CR6_2 Vbiasn1 Vbiasn2 Vbiasp
*.PININFO Vbiasn1:O Vbiasn2:O Vbiasp:O
MM2 Vbiasp Vbiasn2 Vbiasn1 gnd! nmos w=WA l=LA nfin=nA1
MM0 Vbiasn2 Vbiasn1 gnd! gnd! nmos w=WA l=LA nfin=nA2
MM4 Vbiasn1 net15 gnd! gnd! nmos w=WA l=LA nfin=nA3
MM5 net15 net15 gnd! gnd! nmos w=WA l=LA nfin=nA3
MM3 Vbiasp Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA4
MM1 Vbiasn2 Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA4
MM6 net15 Vbiasp vdd! vdd! pmos w=WA l=LA nfin=nA5
.ENDS


xiota LG_Vbiasn1 LG_Vbiasn2 LG_Vbiasp LG_Vbiasp1 LG_Vbiasp2 Vinn Vinp Voutn Voutp fully_differential_folded_cascode_pmos
xiLG_load_biasn_LV LG_Vbiasn2 Biasp LG_load_biasn_LV
xibCR6_2 Biasn1 Biasn2 Biasp CR6_2
.END