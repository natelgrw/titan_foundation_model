.suckt  two_stage_single_output_op_amp_94_4 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorNmos2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorNmos7 out inputVoltageBiasXXnXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mNormalTransistorNmos8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mNormalTransistorNmos9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 sourceTransconductance outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
mNormalTransistorNmos11 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mNormalTransistorNmos12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
mNormalTransistorNmos14 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
mNormalTransistorPmos15 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos16 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos17 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mNormalTransistorPmos18 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mNormalTransistorPmos19 outVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos20 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos
mNormalTransistorPmos21 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_94_4

