.suckt  two_stage_single_output_op_amp_139_12 ibias in1 in2 out sourceNmos sourcePmos
mDiodeTransistorNmos1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mDiodeTransistorNmos2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mDiodeTransistorNmos3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mDiodeTransistorPmos4 ibias ibias sourcePmos sourcePmos pmos
mDiodeTransistorPmos5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mDiodeTransistorPmos6 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mNormalTransistorNmos7 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos8 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mNormalTransistorNmos9 outFirstStage outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos10 FirstStageYinnerOutputLoad1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mNormalTransistorNmos11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mNormalTransistorPmos12 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mNormalTransistorPmos13 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mNormalTransistorPmos14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos15 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos16 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos17 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerOutputLoad1 sourcePmos sourcePmos pmos
mNormalTransistorPmos18 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerOutputLoad1 sourcePmos sourcePmos pmos
mNormalTransistorPmos19 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mNormalTransistorPmos20 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mNormalTransistorPmos21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
Capacitor1 out sourceNmos 
Capacitor2 outFirstStage out 
.end two_stage_single_output_op_amp_139_12

